../../rtl/prim_clock_gating.v